// Copyright (c) 2020 ETH Zurich and University of Bologna
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

import axi_pkg::*;
import pulp_cluster_cfg_pkg::*;

// Stub of PULP Cluster for out-of-context synthesis
module pulp_cluster_ooc (
  input  logic          clk_i,
  input  logic          rst_ni,
  input  logic          ref_clk_i,
  input  cluster_id_t   cluster_id_i,
  input  logic          fetch_en_i,
  output logic          eoc_o,
  output logic          busy_o,

  // Slave Port
  // AW
  input  pulp_cluster_cfg_pkg::addr_t         slv_aw_addr_i,
  input  prot_t         slv_aw_prot_i,
  input  region_t       slv_aw_region_i,
  input  len_t          slv_aw_len_i,
  input  size_t         slv_aw_size_i,
  input  burst_t        slv_aw_burst_i,
  input  logic          slv_aw_lock_i,
  input  atop_t         slv_aw_atop_i,
  input  cache_t        slv_aw_cache_i,
  input  qos_t          slv_aw_qos_i,
  input  id_slv_t       slv_aw_id_i,
  input  pulp_cluster_cfg_pkg::user_t         slv_aw_user_i,
  // used if ASYNC_INTF
  input  dc_buf_t       slv_aw_writetoken_i,
  output dc_buf_t       slv_aw_readpointer_o,
  // used if !ASYNC_INTF
  input  logic          slv_aw_valid_i,
  output logic          slv_aw_ready_o,
  // AR
  input  pulp_cluster_cfg_pkg::addr_t         slv_ar_addr_i,
  input  prot_t         slv_ar_prot_i,
  input  region_t       slv_ar_region_i,
  input  len_t          slv_ar_len_i,
  input  size_t         slv_ar_size_i,
  input  burst_t        slv_ar_burst_i,
  input  logic          slv_ar_lock_i,
  input  cache_t        slv_ar_cache_i,
  input  qos_t          slv_ar_qos_i,
  input  id_slv_t       slv_ar_id_i,
  input  pulp_cluster_cfg_pkg::user_t         slv_ar_user_i,
  // used if ASYNC_INTF
  input  dc_buf_t       slv_ar_writetoken_i,
  output dc_buf_t       slv_ar_readpointer_o,
  // used if !ASYNC_INTF
  input  logic          slv_ar_valid_i,
  output logic          slv_ar_ready_o,
  // W
  input  pulp_cluster_cfg_pkg::data_t         slv_w_data_i,
  input  pulp_cluster_cfg_pkg::strb_t         slv_w_strb_i,
  input  pulp_cluster_cfg_pkg::user_t         slv_w_user_i,
  input  logic          slv_w_last_i,
  // used if ASYNC_INTF
  input  dc_buf_t       slv_w_writetoken_i,
  output dc_buf_t       slv_w_readpointer_o,
  // used if !ASYNC_INTF
  input  logic          slv_w_valid_i,
  output logic          slv_w_ready_o,
  // R
  output pulp_cluster_cfg_pkg::data_t         slv_r_data_o,
  output axi_pkg::resp_t         slv_r_resp_o,
  output logic          slv_r_last_o,
  output id_slv_t       slv_r_id_o,
  output pulp_cluster_cfg_pkg::user_t         slv_r_user_o,
  // used if ASYNC_INTF
  output dc_buf_t       slv_r_writetoken_o,
  input  dc_buf_t       slv_r_readpointer_i,
  // used if !ASYNC_INTF
  output logic          slv_r_valid_o,
  input  logic          slv_r_ready_i,
  // B
  output axi_pkg::resp_t         slv_b_resp_o,
  output id_slv_t       slv_b_id_o,
  output pulp_cluster_cfg_pkg::user_t         slv_b_user_o,
  // used if ASYNC_INTF
  output dc_buf_t       slv_b_writetoken_o,
  input  dc_buf_t       slv_b_readpointer_i,
  // used if !ASYNC_INTF
  output logic          slv_b_valid_o,
  input  logic          slv_b_ready_i,

  // Master Port
  // AW
  output pulp_cluster_cfg_pkg::addr_t         mst_aw_addr_o,
  output prot_t         mst_aw_prot_o,
  output region_t       mst_aw_region_o,
  output len_t          mst_aw_len_o,
  output size_t         mst_aw_size_o,
  output burst_t        mst_aw_burst_o,
  output logic          mst_aw_lock_o,
  output atop_t         mst_aw_atop_o,
  output cache_t        mst_aw_cache_o,
  output qos_t          mst_aw_qos_o,
  output id_mst_t       mst_aw_id_o,
  output pulp_cluster_cfg_pkg::user_t         mst_aw_user_o,
  // used if ASYNC_INTF
  output dc_buf_t       mst_aw_writetoken_o,
  input  dc_buf_t       mst_aw_readpointer_i,
  // used if !ASYNC_INTF
  output logic          mst_aw_valid_o,
  input  logic          mst_aw_ready_i,
  // AR
  output pulp_cluster_cfg_pkg::addr_t         mst_ar_addr_o,
  output prot_t         mst_ar_prot_o,
  output region_t       mst_ar_region_o,
  output len_t          mst_ar_len_o,
  output size_t         mst_ar_size_o,
  output burst_t        mst_ar_burst_o,
  output logic          mst_ar_lock_o,
  output cache_t        mst_ar_cache_o,
  output qos_t          mst_ar_qos_o,
  output id_mst_t       mst_ar_id_o,
  output pulp_cluster_cfg_pkg::user_t         mst_ar_user_o,
  // used if ASYNC_INTF
  output dc_buf_t       mst_ar_writetoken_o,
  input  dc_buf_t       mst_ar_readpointer_i,
  // used if !ASYNC_INTF
  output logic          mst_ar_valid_o,
  input  logic          mst_ar_ready_i,
  // W
  output pulp_cluster_cfg_pkg::data_t         mst_w_data_o,
  output pulp_cluster_cfg_pkg::strb_t         mst_w_strb_o,
  output pulp_cluster_cfg_pkg::user_t         mst_w_user_o,
  output logic          mst_w_last_o,
  // used if ASYNC_INTF
  output dc_buf_t       mst_w_writetoken_o,
  input  dc_buf_t       mst_w_readpointer_i,
  // used if !ASYNC_INTF
  output logic          mst_w_valid_o,
  input  logic          mst_w_ready_i,
  // R
  input  pulp_cluster_cfg_pkg::data_t         mst_r_data_i,
  input  axi_pkg::resp_t         mst_r_resp_i,
  input  logic          mst_r_last_i,
  input  id_mst_t       mst_r_id_i,
  input  pulp_cluster_cfg_pkg::user_t         mst_r_user_i,
  // used if ASYNC_INTF
  input  dc_buf_t       mst_r_writetoken_i,
  output dc_buf_t       mst_r_readpointer_o,
  // used if !ASYNC_INTF
  input  logic          mst_r_valid_i,
  output logic          mst_r_ready_o,
  // B
  input  axi_pkg::resp_t         mst_b_resp_i,
  input  id_mst_t       mst_b_id_i,
  input  pulp_cluster_cfg_pkg::user_t         mst_b_user_i,
  // used if ASYNC_INTF
  input  dc_buf_t       mst_b_writetoken_i,
  output dc_buf_t       mst_b_readpointer_o,
  // used if !ASYNC_INTF
  input  logic          mst_b_valid_i,
  output logic          mst_b_ready_o,

  // AXI4 DMA MASTER
  // WRITE ADDRESS CHANNEL
  output pulp_cluster_cfg_pkg::addr_t         dma_aw_addr_o,
  output prot_t         dma_aw_prot_o,
  output region_t       dma_aw_region_o,
  output len_t          dma_aw_len_o,
  output size_t         dma_aw_size_o,
  output burst_t        dma_aw_burst_o,
  output logic          dma_aw_lock_o,
  output atop_t         dma_aw_atop_o,
  output cache_t        dma_aw_cache_o,
  output qos_t          dma_aw_qos_o,
  output id_dma_t       dma_aw_id_o,
  output pulp_cluster_cfg_pkg::user_t         dma_aw_user_o,
  output logic          dma_aw_valid_o,
  input  logic          dma_aw_ready_i,

  // READ ADDRESS CHANNEL
  output pulp_cluster_cfg_pkg::addr_t         dma_ar_addr_o,
  output prot_t         dma_ar_prot_o,
  output region_t       dma_ar_region_o,
  output len_t          dma_ar_len_o,
  output size_t         dma_ar_size_o,
  output burst_t        dma_ar_burst_o,
  output logic          dma_ar_lock_o,
  output cache_t        dma_ar_cache_o,
  output qos_t          dma_ar_qos_o,
  output id_dma_t       dma_ar_id_o,
  output pulp_cluster_cfg_pkg::user_t         dma_ar_user_o,
  output logic          dma_ar_valid_o,
  input  logic          dma_ar_ready_i,

  // WRITE DATA CHANNEL
  output data_dma_t     dma_w_data_o,
  output strb_dma_t     dma_w_strb_o,
  output pulp_cluster_cfg_pkg::user_t         dma_w_user_o,
  output logic          dma_w_last_o,
  output logic          dma_w_valid_o,
  input  logic          dma_w_ready_i,

  // READ DATA CHANNEL
  input  data_dma_t     dma_r_data_i,
  input  axi_pkg::resp_t         dma_r_resp_i,
  input  logic          dma_r_last_i,
  input  id_dma_t       dma_r_id_i,
  input  pulp_cluster_cfg_pkg::user_t         dma_r_user_i,
  input  logic          dma_r_valid_i,
  output logic          dma_r_ready_o,

  // WRITE RESPONSE CHANNEL
  input  axi_pkg::resp_t         dma_b_resp_i,
  input  id_dma_t       dma_b_id_i,
  input  pulp_cluster_cfg_pkg::user_t         dma_b_user_i,
  input  logic          dma_b_valid_i,
  output logic          dma_b_ready_o,

  //AXI4 NHI SLAVE
  // WRITE ADDRESS CHANNEL
  input  pulp_cluster_cfg_pkg::addr_t         nhi_aw_addr_i,
  input  prot_t         nhi_aw_prot_i,
  input  region_t       nhi_aw_region_i,
  input  len_t          nhi_aw_len_i,
  input  size_t         nhi_aw_size_i,
  input  burst_t        nhi_aw_burst_i,
  input  logic          nhi_aw_lock_i,
  input  atop_t         nhi_aw_atop_i,
  input  cache_t        nhi_aw_cache_i,
  input  qos_t          nhi_aw_qos_i,
  input  id_dma_t       nhi_aw_id_i,
  input  pulp_cluster_cfg_pkg::user_t         nhi_aw_user_i,
  input  logic          nhi_aw_valid_i,
  output logic          nhi_aw_ready_o,

  // READ ADDRESS CHANNEL
  input  pulp_cluster_cfg_pkg::addr_t         nhi_ar_addr_i,
  input  prot_t         nhi_ar_prot_i,
  input  region_t       nhi_ar_region_i,
  input  len_t          nhi_ar_len_i,
  input  size_t         nhi_ar_size_i,
  input  burst_t        nhi_ar_burst_i,
  input  logic          nhi_ar_lock_i,
  input  cache_t        nhi_ar_cache_i,
  input  qos_t          nhi_ar_qos_i,
  input  id_dma_t       nhi_ar_id_i,
  input  pulp_cluster_cfg_pkg::user_t         nhi_ar_user_i,
  input  logic          nhi_ar_valid_i,
  output logic          nhi_ar_ready_o,

  // WRITE DATA CHANNEL
  input  data_dma_t     nhi_w_data_i,
  input  strb_dma_t     nhi_w_strb_i,
  input  pulp_cluster_cfg_pkg::user_t         nhi_w_user_i,
  input  logic          nhi_w_last_i,
  input  logic          nhi_w_valid_i,
  output logic          nhi_w_ready_o,

  // READ DATA CHANNEL
  output data_dma_t     nhi_r_data_o,
  output axi_pkg::resp_t         nhi_r_resp_o,
  output logic          nhi_r_last_o,
  output id_dma_t       nhi_r_id_o,
  output pulp_cluster_cfg_pkg::user_t         nhi_r_user_o,
  output logic          nhi_r_valid_o,
  input  logic          nhi_r_ready_i,

  // WRITE RESPONSE CHANNEL
  output axi_pkg::resp_t         nhi_b_resp_o,
  output id_dma_t       nhi_b_id_o,
  output pulp_cluster_cfg_pkg::user_t         nhi_b_user_o,
  output logic          nhi_b_valid_o,
  input  logic          nhi_b_ready_i,

  // Instruction Cache Master Port
  output pulp_cluster_cfg_pkg::addr_t         icache_aw_addr_o,
  output prot_t         icache_aw_prot_o,
  output region_t       icache_aw_region_o,
  output len_t          icache_aw_len_o,
  output size_t         icache_aw_size_o,
  output burst_t        icache_aw_burst_o,
  output logic          icache_aw_lock_o,
  output atop_t         icache_aw_atop_o,
  output cache_t        icache_aw_cache_o,
  output qos_t          icache_aw_qos_o,
  output id_icache_t    icache_aw_id_o,
  output pulp_cluster_cfg_pkg::user_t         icache_aw_user_o,
  output logic          icache_aw_valid_o,
  input  logic          icache_aw_ready_i,

  output pulp_cluster_cfg_pkg::addr_t         icache_ar_addr_o,
  output prot_t         icache_ar_prot_o,
  output region_t       icache_ar_region_o,
  output len_t          icache_ar_len_o,
  output size_t         icache_ar_size_o,
  output burst_t        icache_ar_burst_o,
  output logic          icache_ar_lock_o,
  output cache_t        icache_ar_cache_o,
  output qos_t          icache_ar_qos_o,
  output id_icache_t    icache_ar_id_o,
  output pulp_cluster_cfg_pkg::user_t         icache_ar_user_o,
  output logic          icache_ar_valid_o,
  input  logic          icache_ar_ready_i,

  output data_icache_t  icache_w_data_o,
  output strb_icache_t  icache_w_strb_o,
  output pulp_cluster_cfg_pkg::user_t         icache_w_user_o,
  output logic          icache_w_last_o,
  output logic          icache_w_valid_o,
  input  logic          icache_w_ready_i,

  input  data_icache_t  icache_r_data_i,
  input  axi_pkg::resp_t         icache_r_resp_i,
  input  logic          icache_r_last_i,
  input  id_icache_t    icache_r_id_i,
  input  pulp_cluster_cfg_pkg::user_t         icache_r_user_i,
  input  logic          icache_r_valid_i,
  output logic          icache_r_ready_o,

  input  axi_pkg::resp_t         icache_b_resp_i,
  input  id_icache_t    icache_b_id_i,
  input  pulp_cluster_cfg_pkg::user_t         icache_b_user_i,
  input  logic          icache_b_valid_i,
  output logic          icache_b_ready_o,

  input  logic                       task_valid_i,
  output logic                       task_ready_o,
  input  pspin_cfg_pkg::handler_task_t   task_descr_i,

  output logic                       feedback_valid_o,
  input  logic                       feedback_ready_i,
  output pspin_cfg_pkg::feedback_descr_t feedback_o,

  output logic                       cluster_active_o,

  input  logic                       cmd_ready_i,
  output logic                       cmd_valid_o,
  output pspin_cfg_pkg::pspin_cmd_t      cmd_o,

  input  logic                       cmd_resp_valid_i,
  input  pspin_cfg_pkg::pspin_cmd_resp_t cmd_resp_i
);

  pulp_cluster #(
    .ASYNC_INTF               (ASYNC),
    .NB_CORES                 (N_CORES),
    .NB_HWACC_PORTS           (0),
    .NB_DMAS                  (N_DMAS),
    .CLUSTER_ALIAS            (1'b1),
    .CLUSTER_ALIAS_BASE       (12'h1B0),
    .TCDM_SIZE                (TCDM_SIZE),
    .NB_TCDM_BANKS            (N_TCDM_BANKS),
    .XNE_PRESENT              (1'b0),
    // I$ Parameters
    .NB_CACHE_BANKS           (4),
    .CACHE_SIZE               (ICACHE_SIZE),
    .L2_SIZE                  (L2_SIZE),
    // Core Parameters
    .DEM_PER_BEFORE_TCDM_TS   (1'b0),
    .ROM_BOOT_ADDR            (32'h1A00_0000),
    .BOOT_ADDR                (32'h1D00_0080),
    // AXI Parameters
    .AXI_ADDR_WIDTH           (AXI_AW),
    .AXI_DATA_C2S_WIDTH       (AXI_DW),
    .AXI_DATA_S2C_WIDTH       (AXI_DW),
    .AXI_USER_WIDTH           (AXI_UW),
    .AXI_ID_IN_WIDTH          (AXI_IW_SLV),
    .AXI_ID_OUT_WIDTH         (AXI_IW_MST),
    .DC_SLICE_BUFFER_WIDTH    (DC_BUF_W),
    // TCDM and Interconnect Parameters
    .DATA_WIDTH               (32),
    .ADDR_WIDTH               (32),
    .TEST_SET_BIT             (20),
    // DMA Parameters
    .NB_OUTSND_BURSTS         (DMA_MAX_N_TXNS),
    .MCHAN_BURST_LENGTH       (DMA_MAX_BURST_SIZE)
  ) i_bound (
    .clk_i,
    .rst_ni,
    .ref_clk_i,

    .pmu_mem_pwdn_i               (1'b0),
    .base_addr_i                  ('0),
    .test_mode_i                  ('0),
    .en_sa_boot_i                 ('0),

    .cluster_id_i,

    .fetch_en_i,
    .eoc_o,
    .busy_o,

    .ext_events_writetoken_i      ('0),
    .ext_events_readpointer_o     (),
    .ext_events_dataasync_i       ('0),
    .dma_pe_evt_ack_i             ('0),
    .dma_pe_evt_valid_o           (),
    .dma_pe_irq_ack_i             ('0),
    .dma_pe_irq_valid_o           (),
    .pf_evt_ack_i                 ('0),
    .pf_evt_valid_o               (),

    .data_slave_aw_addr_i         (slv_aw_addr_i),
    .data_slave_aw_prot_i         (slv_aw_prot_i),
    .data_slave_aw_region_i       (slv_aw_region_i),
    .data_slave_aw_len_i          (slv_aw_len_i),
    .data_slave_aw_size_i         (slv_aw_size_i),
    .data_slave_aw_burst_i        (slv_aw_burst_i),
    .data_slave_aw_lock_i         (slv_aw_lock_i),
    .data_slave_aw_atop_i         (slv_aw_atop_i),
    .data_slave_aw_cache_i        (slv_aw_cache_i),
    .data_slave_aw_qos_i          (slv_aw_qos_i),
    .data_slave_aw_id_i           (slv_aw_id_i),
    .data_slave_aw_user_i         (slv_aw_user_i),
    .data_slave_aw_writetoken_i   (slv_aw_writetoken_i),
    .data_slave_aw_readpointer_o  (slv_aw_readpointer_o),
    .data_slave_aw_valid_i        (slv_aw_valid_i),
    .data_slave_aw_ready_o        (slv_aw_ready_o),
    .data_slave_ar_addr_i         (slv_ar_addr_i),
    .data_slave_ar_prot_i         (slv_ar_prot_i),
    .data_slave_ar_region_i       (slv_ar_region_i),
    .data_slave_ar_len_i          (slv_ar_len_i),
    .data_slave_ar_size_i         (slv_ar_size_i),
    .data_slave_ar_burst_i        (slv_ar_burst_i),
    .data_slave_ar_lock_i         (slv_ar_lock_i),
    .data_slave_ar_cache_i        (slv_ar_cache_i),
    .data_slave_ar_qos_i          (slv_ar_qos_i),
    .data_slave_ar_id_i           (slv_ar_id_i),
    .data_slave_ar_user_i         (slv_ar_user_i),
    .data_slave_ar_writetoken_i   (slv_ar_writetoken_i),
    .data_slave_ar_readpointer_o  (slv_ar_readpointer_o),
    .data_slave_ar_valid_i        (slv_ar_valid_i),
    .data_slave_ar_ready_o        (slv_ar_ready_o),
    .data_slave_w_data_i          (slv_w_data_i),
    .data_slave_w_strb_i          (slv_w_strb_i),
    .data_slave_w_user_i          (slv_w_user_i),
    .data_slave_w_last_i          (slv_w_last_i),
    .data_slave_w_writetoken_i    (slv_w_writetoken_i),
    .data_slave_w_readpointer_o   (slv_w_readpointer_o),
    .data_slave_w_valid_i         (slv_w_valid_i),
    .data_slave_w_ready_o         (slv_w_ready_o),
    .data_slave_r_data_o          (slv_r_data_o),
    .data_slave_r_resp_o          (slv_r_resp_o),
    .data_slave_r_last_o          (slv_r_last_o),
    .data_slave_r_id_o            (slv_r_id_o),
    .data_slave_r_user_o          (slv_r_user_o),
    .data_slave_r_writetoken_o    (slv_r_writetoken_o),
    .data_slave_r_readpointer_i   (slv_r_readpointer_i),
    .data_slave_r_valid_o         (slv_r_valid_o),
    .data_slave_r_ready_i         (slv_r_ready_i),
    .data_slave_b_resp_o          (slv_b_resp_o),
    .data_slave_b_id_o            (slv_b_id_o),
    .data_slave_b_user_o          (slv_b_user_o),
    .data_slave_b_writetoken_o    (slv_b_writetoken_o),
    .data_slave_b_readpointer_i   (slv_b_readpointer_i),
    .data_slave_b_valid_o         (slv_b_valid_o),
    .data_slave_b_ready_i         (slv_b_ready_i),

    .data_master_aw_addr_o        (mst_aw_addr_o),
    .data_master_aw_prot_o        (mst_aw_prot_o),
    .data_master_aw_region_o      (mst_aw_region_o),
    .data_master_aw_len_o         (mst_aw_len_o),
    .data_master_aw_size_o        (mst_aw_size_o),
    .data_master_aw_burst_o       (mst_aw_burst_o),
    .data_master_aw_lock_o        (mst_aw_lock_o),
    .data_master_aw_atop_o        (mst_aw_atop_o),
    .data_master_aw_cache_o       (),
    .data_master_aw_qos_o         (mst_aw_qos_o),
    .data_master_aw_id_o          (mst_aw_id_o),
    .data_master_aw_user_o        (mst_aw_user_o),
    .data_master_aw_writetoken_o  (mst_aw_writetoken_o),
    .data_master_aw_readpointer_i (mst_aw_readpointer_i),
    .data_master_aw_valid_o       (mst_aw_valid_o),
    .data_master_aw_ready_i       (mst_aw_ready_i),
    .data_master_ar_addr_o        (mst_ar_addr_o),
    .data_master_ar_prot_o        (mst_ar_prot_o),
    .data_master_ar_region_o      (mst_ar_region_o),
    .data_master_ar_len_o         (mst_ar_len_o),
    .data_master_ar_size_o        (mst_ar_size_o),
    .data_master_ar_burst_o       (mst_ar_burst_o),
    .data_master_ar_lock_o        (mst_ar_lock_o),
    .data_master_ar_cache_o       (),
    .data_master_ar_qos_o         (mst_ar_qos_o),
    .data_master_ar_id_o          (mst_ar_id_o),
    .data_master_ar_user_o        (mst_ar_user_o),
    .data_master_ar_writetoken_o  (mst_ar_writetoken_o),
    .data_master_ar_readpointer_i (mst_ar_readpointer_i),
    .data_master_ar_valid_o       (mst_ar_valid_o),
    .data_master_ar_ready_i       (mst_ar_ready_i),
    .data_master_w_data_o         (mst_w_data_o),
    .data_master_w_strb_o         (mst_w_strb_o),
    .data_master_w_user_o         (mst_w_user_o),
    .data_master_w_last_o         (mst_w_last_o),
    .data_master_w_writetoken_o   (mst_w_writetoken_o),
    .data_master_w_readpointer_i  (mst_w_readpointer_i),
    .data_master_w_valid_o        (mst_w_valid_o),
    .data_master_w_ready_i        (mst_w_ready_i),
    .data_master_r_data_i         (mst_r_data_i),
    .data_master_r_resp_i         (mst_r_resp_i),
    .data_master_r_last_i         (mst_r_last_i),
    .data_master_r_id_i           (mst_r_id_i),
    .data_master_r_user_i         (mst_r_user_i),
    .data_master_r_writetoken_i   (mst_r_writetoken_i),
    .data_master_r_readpointer_o  (mst_r_readpointer_o),
    .data_master_r_valid_i        (mst_r_valid_i),
    .data_master_r_ready_o        (mst_r_ready_o),
    .data_master_b_resp_i         (mst_b_resp_i),
    .data_master_b_id_i           (mst_b_id_i),
    .data_master_b_user_i         (mst_b_user_i),
    .data_master_b_writetoken_i   (mst_b_writetoken_i),
    .data_master_b_readpointer_o  (mst_b_readpointer_o),
    .data_master_b_valid_i        (mst_b_valid_i),
    .data_master_b_ready_o        (mst_b_ready_o),

    .dma_aw_addr_o,
    .dma_aw_prot_o,
    .dma_aw_region_o,
    .dma_aw_len_o,
    .dma_aw_size_o,
    .dma_aw_burst_o,
    .dma_aw_lock_o,
    .dma_aw_atop_o,
    .dma_aw_cache_o   (),
    .dma_aw_qos_o,
    .dma_aw_id_o,
    .dma_aw_user_o,
    .dma_aw_valid_o,
    .dma_aw_ready_i,
    .dma_ar_addr_o,
    .dma_ar_prot_o,
    .dma_ar_region_o,
    .dma_ar_len_o,
    .dma_ar_size_o,
    .dma_ar_burst_o,
    .dma_ar_lock_o,
    .dma_ar_cache_o   (),
    .dma_ar_qos_o,
    .dma_ar_id_o,
    .dma_ar_user_o,
    .dma_ar_valid_o,
    .dma_ar_ready_i,
    .dma_w_data_o,
    .dma_w_strb_o,
    .dma_w_user_o,
    .dma_w_last_o,
    .dma_w_valid_o,
    .dma_w_ready_i,
    .dma_r_data_i,
    .dma_r_resp_i,
    .dma_r_last_i,
    .dma_r_id_i,
    .dma_r_user_i,
    .dma_r_valid_i,
    .dma_r_ready_o,
    .dma_b_resp_i,
    .dma_b_id_i,
    .dma_b_user_i,
    .dma_b_valid_i,
    .dma_b_ready_o,

    .nhi_aw_addr_i,
    .nhi_aw_prot_i,
    .nhi_aw_region_i,
    .nhi_aw_len_i,
    .nhi_aw_size_i,
    .nhi_aw_burst_i,
    .nhi_aw_lock_i,
    .nhi_aw_atop_i,
    .nhi_aw_cache_i,
    .nhi_aw_qos_i,
    .nhi_aw_id_i,
    .nhi_aw_user_i,
    .nhi_aw_valid_i,
    .nhi_aw_ready_o,
    .nhi_ar_addr_i,
    .nhi_ar_prot_i,
    .nhi_ar_region_i,
    .nhi_ar_len_i,
    .nhi_ar_size_i,
    .nhi_ar_burst_i,
    .nhi_ar_lock_i,
    .nhi_ar_cache_i,
    .nhi_ar_qos_i,
    .nhi_ar_id_i,
    .nhi_ar_user_i,
    .nhi_ar_valid_i,
    .nhi_ar_ready_o,
    .nhi_w_data_i,
    .nhi_w_strb_i,
    .nhi_w_user_i,
    .nhi_w_last_i,
    .nhi_w_valid_i,
    .nhi_w_ready_o,
    .nhi_r_data_o,
    .nhi_r_resp_o,
    .nhi_r_last_o,
    .nhi_r_id_o,
    .nhi_r_user_o,
    .nhi_r_valid_o,
    .nhi_r_ready_i,
    .nhi_b_resp_o,
    .nhi_b_id_o,
    .nhi_b_user_o,
    .nhi_b_valid_o,
    .nhi_b_ready_i,

    .icache_aw_addr_o,
    .icache_aw_prot_o,
    .icache_aw_region_o,
    .icache_aw_len_o,
    .icache_aw_size_o,
    .icache_aw_burst_o,
    .icache_aw_lock_o,
    .icache_aw_atop_o,
    .icache_aw_cache_o,
    .icache_aw_qos_o,
    .icache_aw_id_o,
    .icache_aw_user_o,
    .icache_aw_valid_o,
    .icache_aw_ready_i,
    .icache_ar_addr_o,
    .icache_ar_prot_o,
    .icache_ar_region_o,
    .icache_ar_len_o,
    .icache_ar_size_o,
    .icache_ar_burst_o,
    .icache_ar_lock_o,
    .icache_ar_cache_o,
    .icache_ar_qos_o,
    .icache_ar_id_o,
    .icache_ar_user_o,
    .icache_ar_valid_o,
    .icache_ar_ready_i,
    .icache_w_data_o,
    .icache_w_strb_o,
    .icache_w_user_o,
    .icache_w_last_o,
    .icache_w_valid_o,
    .icache_w_ready_i,
    .icache_r_data_i,
    .icache_r_resp_i,
    .icache_r_last_i,
    .icache_r_id_i,
    .icache_r_user_i,
    .icache_r_valid_i,
    .icache_r_ready_o,
    .icache_b_resp_i,
    .icache_b_id_i,
    .icache_b_user_i,
    .icache_b_valid_i,
    .icache_b_ready_o,

    .task_valid_i         (task_valid_i),
    .task_ready_o         (task_ready_o),
    .task_descr_i         (task_descr_i),
    .feedback_valid_o     (feedback_valid_o),
    .feedback_ready_i     (feedback_ready_i),
    .feedback_o           (feedback_o),
    .cluster_active_o     (cluster_active_o),
    .cmd_ready_i          (cmd_ready_i),
    .cmd_valid_o          (cmd_valid_o),
    .cmd_o                (cmd_o),
    .cmd_resp_valid_i     (cmd_resp_valid_i),
    .cmd_resp_i           (cmd_resp_i)
  );
  // Make all reads and writes from cluster modifiable.
  // TODO: This might be undesired for transactions from cores to peripherals, better modify the
  // DMA and I$ to issue modifiable transactions.
  assign mst_ar_cache_o = 4'b0010;
  assign mst_aw_cache_o = 4'b0010;
  assign dma_ar_cache_o = 4'b0010;
  assign dma_aw_cache_o = 4'b0010;

endmodule


// Interface wrapper for OOC-synthesized synchronous PULP cluster
module pulp_cluster_sync (
  input  logic        clk_i,
  input  logic        rst_ni,
  input  logic        ref_clk_i,
  input  cluster_id_t cluster_id_i,
  input  logic        fetch_en_i,
  output logic        eoc_o,
  output logic        busy_o,
  AXI_BUS.Slave       slv,
  AXI_BUS.Master      mst,
  AXI_BUS.Master      dma,
  AXI_BUS.Master      icache,
  AXI_BUS.Slave       nhi,

  input  logic                       task_valid_i,
  output logic                       task_ready_o,
  input  pspin_cfg_pkg::handler_task_t   task_descr_i,
  output logic                       feedback_valid_o,
  input  logic                       feedback_ready_i,
  output pspin_cfg_pkg::feedback_descr_t feedback_o,
  output logic                       cluster_active_o,
  input  logic                       cmd_ready_i,
  output logic                       cmd_valid_o,
  output pspin_cfg_pkg::pspin_cmd_t      cmd_o,
  input  logic                       cmd_resp_valid_i,
  input  pspin_cfg_pkg::pspin_cmd_resp_t cmd_resp_i
);

  pulp_cluster_ooc i_ooc (
    .clk_i,
    .rst_ni,
    .ref_clk_i,
    .cluster_id_i,
    .fetch_en_i,
    .eoc_o,
    .busy_o,

    .slv_aw_addr_i        (slv.aw_addr),
    .slv_aw_prot_i        (slv.aw_prot),
    .slv_aw_region_i      (slv.aw_region),
    .slv_aw_len_i         (slv.aw_len),
    .slv_aw_size_i        (slv.aw_size),
    .slv_aw_burst_i       (slv.aw_burst),
    .slv_aw_lock_i        (slv.aw_lock),
    .slv_aw_atop_i        (slv.aw_atop),
    .slv_aw_cache_i       (slv.aw_cache),
    .slv_aw_qos_i         (slv.aw_qos),
    .slv_aw_id_i          (slv.aw_id),
    .slv_aw_user_i        (slv.aw_user),
    .slv_aw_valid_i       (slv.aw_valid),
    .slv_aw_ready_o       (slv.aw_ready),
    .slv_aw_writetoken_i  (),
    .slv_aw_readpointer_o (),
    .slv_ar_addr_i        (slv.ar_addr),
    .slv_ar_prot_i        (slv.ar_prot),
    .slv_ar_region_i      (slv.ar_region),
    .slv_ar_len_i         (slv.ar_len),
    .slv_ar_size_i        (slv.ar_size),
    .slv_ar_burst_i       (slv.ar_burst),
    .slv_ar_lock_i        (slv.ar_lock),
    .slv_ar_cache_i       (slv.ar_cache),
    .slv_ar_qos_i         (slv.ar_qos),
    .slv_ar_id_i          (slv.ar_id),
    .slv_ar_user_i        (slv.ar_user),
    .slv_ar_valid_i       (slv.ar_valid),
    .slv_ar_ready_o       (slv.ar_ready),
    .slv_ar_writetoken_i  (),
    .slv_ar_readpointer_o (),
    .slv_w_data_i         (slv.w_data),
    .slv_w_strb_i         (slv.w_strb),
    .slv_w_user_i         (slv.w_user),
    .slv_w_last_i         (slv.w_last),
    .slv_w_valid_i        (slv.w_valid),
    .slv_w_ready_o        (slv.w_ready),
    .slv_w_writetoken_i   (),
    .slv_w_readpointer_o  (),
    .slv_r_data_o         (slv.r_data),
    .slv_r_resp_o         (slv.r_resp),
    .slv_r_last_o         (slv.r_last),
    .slv_r_id_o           (slv.r_id),
    .slv_r_user_o         (slv.r_user),
    .slv_r_valid_o        (slv.r_valid),
    .slv_r_ready_i        (slv.r_ready),
    .slv_r_writetoken_o   (),
    .slv_r_readpointer_i  (),
    .slv_b_resp_o         (slv.b_resp),
    .slv_b_id_o           (slv.b_id),
    .slv_b_user_o         (slv.b_user),
    .slv_b_valid_o        (slv.b_valid),
    .slv_b_ready_i        (slv.b_ready),
    .slv_b_writetoken_o   (),
    .slv_b_readpointer_i  (),

    .mst_aw_addr_o        (mst.aw_addr),
    .mst_aw_prot_o        (mst.aw_prot),
    .mst_aw_region_o      (mst.aw_region),
    .mst_aw_len_o         (mst.aw_len),
    .mst_aw_size_o        (mst.aw_size),
    .mst_aw_burst_o       (mst.aw_burst),
    .mst_aw_lock_o        (mst.aw_lock),
    .mst_aw_atop_o        (mst.aw_atop),
    .mst_aw_cache_o       (mst.aw_cache),
    .mst_aw_qos_o         (mst.aw_qos),
    .mst_aw_id_o          (mst.aw_id),
    .mst_aw_user_o        (mst.aw_user),
    .mst_aw_valid_o       (mst.aw_valid),
    .mst_aw_ready_i       (mst.aw_ready),
    .mst_aw_writetoken_o  (),
    .mst_aw_readpointer_i (),
    .mst_ar_addr_o        (mst.ar_addr),
    .mst_ar_prot_o        (mst.ar_prot),
    .mst_ar_region_o      (mst.ar_region),
    .mst_ar_len_o         (mst.ar_len),
    .mst_ar_size_o        (mst.ar_size),
    .mst_ar_burst_o       (mst.ar_burst),
    .mst_ar_lock_o        (mst.ar_lock),
    .mst_ar_cache_o       (mst.ar_cache),
    .mst_ar_qos_o         (mst.ar_qos),
    .mst_ar_id_o          (mst.ar_id),
    .mst_ar_user_o        (mst.ar_user),
    .mst_ar_valid_o       (mst.ar_valid),
    .mst_ar_ready_i       (mst.ar_ready),
    .mst_ar_writetoken_o  (),
    .mst_ar_readpointer_i (),
    .mst_w_data_o         (mst.w_data),
    .mst_w_strb_o         (mst.w_strb),
    .mst_w_user_o         (mst.w_user),
    .mst_w_last_o         (mst.w_last),
    .mst_w_valid_o        (mst.w_valid),
    .mst_w_ready_i        (mst.w_ready),
    .mst_w_writetoken_o   (),
    .mst_w_readpointer_i  (),
    .mst_r_data_i         (mst.r_data),
    .mst_r_resp_i         (mst.r_resp),
    .mst_r_last_i         (mst.r_last),
    .mst_r_id_i           (mst.r_id),
    .mst_r_user_i         (mst.r_user),
    .mst_r_valid_i        (mst.r_valid),
    .mst_r_ready_o        (mst.r_ready),
    .mst_r_writetoken_i   (),
    .mst_r_readpointer_o  (),
    .mst_b_resp_i         (mst.b_resp),
    .mst_b_id_i           (mst.b_id),
    .mst_b_user_i         (mst.b_user),
    .mst_b_valid_i        (mst.b_valid),
    .mst_b_ready_o        (mst.b_ready),
    .mst_b_writetoken_i   (),
    .mst_b_readpointer_o  (),

    .dma_aw_addr_o   (dma.aw_addr),
    .dma_aw_prot_o   (dma.aw_prot),
    .dma_aw_region_o (dma.aw_region),
    .dma_aw_len_o    (dma.aw_len),
    .dma_aw_size_o   (dma.aw_size),
    .dma_aw_burst_o  (dma.aw_burst),
    .dma_aw_lock_o   (dma.aw_lock),
    .dma_aw_atop_o   (dma.aw_atop),
    .dma_aw_cache_o  (dma.aw_cache),
    .dma_aw_qos_o    (dma.aw_qos),
    .dma_aw_id_o     (dma.aw_id),
    .dma_aw_user_o   (dma.aw_user),
    .dma_aw_valid_o  (dma.aw_valid),
    .dma_aw_ready_i  (dma.aw_ready),
    .dma_ar_addr_o   (dma.ar_addr),
    .dma_ar_prot_o   (dma.ar_prot),
    .dma_ar_region_o (dma.ar_region),
    .dma_ar_len_o    (dma.ar_len),
    .dma_ar_size_o   (dma.ar_size),
    .dma_ar_burst_o  (dma.ar_burst),
    .dma_ar_lock_o   (dma.ar_lock),
    .dma_ar_cache_o  (dma.ar_cache),
    .dma_ar_qos_o    (dma.ar_qos),
    .dma_ar_id_o     (dma.ar_id),
    .dma_ar_user_o   (dma.ar_user),
    .dma_ar_valid_o  (dma.ar_valid),
    .dma_ar_ready_i  (dma.ar_ready),
    .dma_w_data_o    (dma.w_data),
    .dma_w_strb_o    (dma.w_strb),
    .dma_w_user_o    (dma.w_user),
    .dma_w_last_o    (dma.w_last),
    .dma_w_valid_o   (dma.w_valid),
    .dma_w_ready_i   (dma.w_ready),
    .dma_r_data_i    (dma.r_data),
    .dma_r_resp_i    (dma.r_resp),
    .dma_r_last_i    (dma.r_last),
    .dma_r_id_i      (dma.r_id),
    .dma_r_user_i    (dma.r_user),
    .dma_r_valid_i   (dma.r_valid),
    .dma_r_ready_o   (dma.r_ready),
    .dma_b_resp_i    (dma.b_resp),
    .dma_b_id_i      (dma.b_id),
    .dma_b_user_i    (dma.b_user),
    .dma_b_valid_i   (dma.b_valid),
    .dma_b_ready_o   (dma.b_ready),

    .nhi_aw_addr_i   (nhi.aw_addr),
    .nhi_aw_prot_i   (nhi.aw_prot),
    .nhi_aw_region_i (nhi.aw_region),
    .nhi_aw_len_i    (nhi.aw_len),
    .nhi_aw_size_i   (nhi.aw_size),
    .nhi_aw_burst_i  (nhi.aw_burst),
    .nhi_aw_lock_i   (nhi.aw_lock),
    .nhi_aw_atop_i   (nhi.aw_atop),
    .nhi_aw_cache_i  (nhi.aw_cache),
    .nhi_aw_qos_i    (nhi.aw_qos),
    .nhi_aw_id_i     (nhi.aw_id),
    .nhi_aw_user_i   (nhi.aw_user),
    .nhi_aw_valid_i  (nhi.aw_valid),
    .nhi_aw_ready_o  (nhi.aw_ready),
    .nhi_ar_addr_i   (nhi.ar_addr),
    .nhi_ar_prot_i   (nhi.ar_prot),
    .nhi_ar_region_i (nhi.ar_region),
    .nhi_ar_len_i    (nhi.ar_len),
    .nhi_ar_size_i   (nhi.ar_size),
    .nhi_ar_burst_i  (nhi.ar_burst),
    .nhi_ar_lock_i   (nhi.ar_lock),
    .nhi_ar_cache_i  (nhi.ar_cache),
    .nhi_ar_qos_i    (nhi.ar_qos),
    .nhi_ar_id_i     (nhi.ar_id),
    .nhi_ar_user_i   (nhi.ar_user),
    .nhi_ar_valid_i  (nhi.ar_valid),
    .nhi_ar_ready_o  (nhi.ar_ready),
    .nhi_w_data_i    (nhi.w_data),
    .nhi_w_strb_i    (nhi.w_strb),
    .nhi_w_user_i    (nhi.w_user),
    .nhi_w_last_i    (nhi.w_last),
    .nhi_w_valid_i   (nhi.w_valid),
    .nhi_w_ready_o   (nhi.w_ready),
    .nhi_r_data_o    (nhi.r_data),
    .nhi_r_resp_o    (nhi.r_resp),
    .nhi_r_last_o    (nhi.r_last),
    .nhi_r_id_o      (nhi.r_id),
    .nhi_r_user_o    (nhi.r_user),
    .nhi_r_valid_o   (nhi.r_valid),
    .nhi_r_ready_i   (nhi.r_ready),
    .nhi_b_resp_o    (nhi.b_resp),
    .nhi_b_id_o      (nhi.b_id),
    .nhi_b_user_o    (nhi.b_user),
    .nhi_b_valid_o   (nhi.b_valid),
    .nhi_b_ready_i   (nhi.b_ready),

    .icache_aw_addr_o   (icache.aw_addr),
    .icache_aw_prot_o   (icache.aw_prot),
    .icache_aw_region_o (icache.aw_region),
    .icache_aw_len_o    (icache.aw_len),
    .icache_aw_size_o   (icache.aw_size),
    .icache_aw_burst_o  (icache.aw_burst),
    .icache_aw_lock_o   (icache.aw_lock),
    .icache_aw_atop_o   (icache.aw_atop),
    .icache_aw_cache_o  (icache.aw_cache),
    .icache_aw_qos_o    (icache.aw_qos),
    .icache_aw_id_o     (icache.aw_id),
    .icache_aw_user_o   (icache.aw_user),
    .icache_aw_valid_o  (icache.aw_valid),
    .icache_aw_ready_i  (icache.aw_ready),
    .icache_ar_addr_o   (icache.ar_addr),
    .icache_ar_prot_o   (icache.ar_prot),
    .icache_ar_region_o (icache.ar_region),
    .icache_ar_len_o    (icache.ar_len),
    .icache_ar_size_o   (icache.ar_size),
    .icache_ar_burst_o  (icache.ar_burst),
    .icache_ar_lock_o   (icache.ar_lock),
    .icache_ar_cache_o  (icache.ar_cache),
    .icache_ar_qos_o    (icache.ar_qos),
    .icache_ar_id_o     (icache.ar_id),
    .icache_ar_user_o   (icache.ar_user),
    .icache_ar_valid_o  (icache.ar_valid),
    .icache_ar_ready_i  (icache.ar_ready),
    .icache_w_data_o    (icache.w_data),
    .icache_w_strb_o    (icache.w_strb),
    .icache_w_user_o    (icache.w_user),
    .icache_w_last_o    (icache.w_last),
    .icache_w_valid_o   (icache.w_valid),
    .icache_w_ready_i   (icache.w_ready),
    .icache_r_data_i    (icache.r_data),
    .icache_r_resp_i    (icache.r_resp),
    .icache_r_last_i    (icache.r_last),
    .icache_r_id_i      (icache.r_id),
    .icache_r_user_i    (icache.r_user),
    .icache_r_valid_i   (icache.r_valid),
    .icache_r_ready_o   (icache.r_ready),
    .icache_b_resp_i    (icache.b_resp),
    .icache_b_id_i      (icache.b_id),
    .icache_b_user_i    (icache.b_user),
    .icache_b_valid_i   (icache.b_valid),
    .icache_b_ready_o   (icache.b_ready),

    .task_valid_i         (task_valid_i),
    .task_ready_o         (task_ready_o),
    .task_descr_i         (task_descr_i),
    .feedback_valid_o     (feedback_valid_o),
    .feedback_ready_i     (feedback_ready_i),
    .feedback_o           (feedback_o),
    .cluster_active_o     (cluster_active_o),
    .cmd_ready_i          (cmd_ready_i),
    .cmd_valid_o          (cmd_valid_o),
    .cmd_o                (cmd_o),
    .cmd_resp_valid_i     (cmd_resp_valid_i),
    .cmd_resp_i           (cmd_resp_i)
  );
endmodule

// Interface wrapper for OOC-synthesized asynchronous PULP cluster
module pulp_cluster_async (
  input  logic          clk_i,
  input  logic          rst_ni,
  input  logic          ref_clk_i,
  input  cluster_id_t   cluster_id_i,
  input  logic          fetch_en_i,
  output logic          eoc_o,
  output logic          busy_o,
  AXI_BUS_ASYNC.Slave   slv,
  AXI_BUS_ASYNC.Master  mst,
  AXI_BUS_ASYNC.Master  dma,
  AXI_BUS_ASYNC.Master  icache
);

  pulp_cluster_ooc i_ooc (
    .clk_i,
    .rst_ni,
    .ref_clk_i,
    .cluster_id_i,
    .fetch_en_i,
    .eoc_o,
    .busy_o,

    .slv_aw_addr_i        (slv.aw_addr),
    .slv_aw_prot_i        (slv.aw_prot),
    .slv_aw_region_i      (slv.aw_region),
    .slv_aw_len_i         (slv.aw_len),
    .slv_aw_size_i        (slv.aw_size),
    .slv_aw_burst_i       (slv.aw_burst),
    .slv_aw_lock_i        (slv.aw_lock),
    .slv_aw_atop_i        (slv.aw_atop),
    .slv_aw_cache_i       (slv.aw_cache),
    .slv_aw_qos_i         (slv.aw_qos),
    .slv_aw_id_i          (slv.aw_id),
    .slv_aw_user_i        (slv.aw_user),
    .slv_aw_valid_i       (),
    .slv_aw_ready_o       (),
    .slv_aw_writetoken_i  (slv.aw_writetoken),
    .slv_aw_readpointer_o (slv.aw_readpointer),
    .slv_ar_addr_i        (slv.ar_addr),
    .slv_ar_prot_i        (slv.ar_prot),
    .slv_ar_region_i      (slv.ar_region),
    .slv_ar_len_i         (slv.ar_len),
    .slv_ar_size_i        (slv.ar_size),
    .slv_ar_burst_i       (slv.ar_burst),
    .slv_ar_lock_i        (slv.ar_lock),
    .slv_ar_cache_i       (slv.ar_cache),
    .slv_ar_qos_i         (slv.ar_qos),
    .slv_ar_id_i          (slv.ar_id),
    .slv_ar_user_i        (slv.ar_user),
    .slv_ar_valid_i       (),
    .slv_ar_ready_o       (),
    .slv_ar_writetoken_i  (slv.ar_writetoken),
    .slv_ar_readpointer_o (slv.ar_readpointer),
    .slv_w_data_i         (slv.w_data),
    .slv_w_strb_i         (slv.w_strb),
    .slv_w_user_i         (slv.w_user),
    .slv_w_last_i         (slv.w_last),
    .slv_w_valid_i        (),
    .slv_w_ready_o        (),
    .slv_w_writetoken_i   (slv.w_writetoken),
    .slv_w_readpointer_o  (slv.w_readpointer),
    .slv_r_data_o         (slv.r_data),
    .slv_r_resp_o         (slv.r_resp),
    .slv_r_last_o         (slv.r_last),
    .slv_r_id_o           (slv.r_id),
    .slv_r_user_o         (slv.r_user),
    .slv_r_valid_o        (),
    .slv_r_ready_i        (),
    .slv_r_writetoken_o   (slv.r_writetoken),
    .slv_r_readpointer_i  (slv.r_readpointer),
    .slv_b_resp_o         (slv.b_resp),
    .slv_b_id_o           (slv.b_id),
    .slv_b_user_o         (slv.b_user),
    .slv_b_valid_o        (),
    .slv_b_ready_i        (),
    .slv_b_writetoken_o   (slv.b_writetoken),
    .slv_b_readpointer_i  (slv.b_readpointer),

    .mst_aw_addr_o        (mst.aw_addr),
    .mst_aw_prot_o        (mst.aw_prot),
    .mst_aw_region_o      (mst.aw_region),
    .mst_aw_len_o         (mst.aw_len),
    .mst_aw_size_o        (mst.aw_size),
    .mst_aw_burst_o       (mst.aw_burst),
    .mst_aw_lock_o        (mst.aw_lock),
    .mst_aw_atop_o        (mst.aw_atop),
    .mst_aw_cache_o       (mst.aw_cache),
    .mst_aw_qos_o         (mst.aw_qos),
    .mst_aw_id_o          (mst.aw_id),
    .mst_aw_user_o        (mst.aw_user),
    .mst_aw_valid_o       (),
    .mst_aw_ready_i       (),
    .mst_aw_writetoken_o  (mst.aw_writetoken),
    .mst_aw_readpointer_i (mst.aw_readpointer),
    .mst_ar_addr_o        (mst.ar_addr),
    .mst_ar_prot_o        (mst.ar_prot),
    .mst_ar_region_o      (mst.ar_region),
    .mst_ar_len_o         (mst.ar_len),
    .mst_ar_size_o        (mst.ar_size),
    .mst_ar_burst_o       (mst.ar_burst),
    .mst_ar_lock_o        (mst.ar_lock),
    .mst_ar_cache_o       (mst.ar_cache),
    .mst_ar_qos_o         (mst.ar_qos),
    .mst_ar_id_o          (mst.ar_id),
    .mst_ar_user_o        (mst.ar_user),
    .mst_ar_valid_o       (),
    .mst_ar_ready_i       (),
    .mst_ar_writetoken_o  (mst.ar_writetoken),
    .mst_ar_readpointer_i (mst.ar_readpointer),
    .mst_w_data_o         (mst.w_data),
    .mst_w_strb_o         (mst.w_strb),
    .mst_w_user_o         (mst.w_user),
    .mst_w_last_o         (mst.w_last),
    .mst_w_valid_o        (),
    .mst_w_ready_i        (),
    .mst_w_writetoken_o   (mst.w_writetoken),
    .mst_w_readpointer_i  (mst.w_readpointer),
    .mst_r_data_i         (mst.r_data),
    .mst_r_resp_i         (mst.r_resp),
    .mst_r_last_i         (mst.r_last),
    .mst_r_id_i           (mst.r_id),
    .mst_r_user_i         (mst.r_user),
    .mst_r_valid_i        (),
    .mst_r_ready_o        (),
    .mst_r_writetoken_i   (mst.r_writetoken),
    .mst_r_readpointer_o  (mst.r_readpointer),
    .mst_b_resp_i         (mst.b_resp),
    .mst_b_id_i           (mst.b_id),
    .mst_b_user_i         (mst.b_user),
    .mst_b_valid_i        (),
    .mst_b_ready_o        (),
    .mst_b_writetoken_i   (mst.b_writetoken),
    .mst_b_readpointer_o  (mst.b_readpointer),

    .dma_aw_addr_o   (dma.aw_addr),
    .dma_aw_prot_o   (dma.aw_prot),
    .dma_aw_region_o (dma.aw_region),
    .dma_aw_len_o    (dma.aw_len),
    .dma_aw_size_o   (dma.aw_size),
    .dma_aw_burst_o  (dma.aw_burst),
    .dma_aw_lock_o   (dma.aw_lock),
    .dma_aw_atop_o   (dma.aw_atop),
    .dma_aw_cache_o  (dma.aw_cache),
    .dma_aw_qos_o    (dma.aw_qos),
    .dma_aw_id_o     (dma.aw_id),
    .dma_aw_user_o   (dma.aw_user),
    .dma_aw_valid_o  (),
    .dma_aw_ready_i  (),
    .dma_ar_addr_o   (dma.ar_addr),
    .dma_ar_prot_o   (dma.ar_prot),
    .dma_ar_region_o (dma.ar_region),
    .dma_ar_len_o    (dma.ar_len),
    .dma_ar_size_o   (dma.ar_size),
    .dma_ar_burst_o  (dma.ar_burst),
    .dma_ar_lock_o   (dma.ar_lock),
    .dma_ar_cache_o  (dma.ar_cache),
    .dma_ar_qos_o    (dma.ar_qos),
    .dma_ar_id_o     (dma.ar_id),
    .dma_ar_user_o   (dma.ar_user),
    .dma_ar_valid_o  (),
    .dma_ar_ready_i  (),
    .dma_w_data_o    (dma.w_data),
    .dma_w_strb_o    (dma.w_strb),
    .dma_w_user_o    (dma.w_user),
    .dma_w_last_o    (dma.w_last),
    .dma_w_valid_o   (),
    .dma_w_ready_i   (),
    .dma_r_data_i    (dma.r_data),
    .dma_r_resp_i    (dma.r_resp),
    .dma_r_last_i    (dma.r_last),
    .dma_r_id_i      (dma.r_id),
    .dma_r_user_i    (dma.r_user),
    .dma_r_valid_i   (),
    .dma_r_ready_o   (),
    .dma_b_resp_i    (dma.b_resp),
    .dma_b_id_i      (dma.b_id),
    .dma_b_user_i    (dma.b_user),
    .dma_b_valid_i   (),
    .dma_b_ready_o   (),

    .icache_aw_addr_o   (icache.aw_addr),
    .icache_aw_prot_o   (icache.aw_prot),
    .icache_aw_region_o (icache.aw_region),
    .icache_aw_len_o    (icache.aw_len),
    .icache_aw_size_o   (icache.aw_size),
    .icache_aw_burst_o  (icache.aw_burst),
    .icache_aw_lock_o   (icache.aw_lock),
    .icache_aw_atop_o   (icache.aw_atop),
    .icache_aw_cache_o  (icache.aw_cache),
    .icache_aw_qos_o    (icache.aw_qos),
    .icache_aw_id_o     (icache.aw_id),
    .icache_aw_user_o   (icache.aw_user),
    .icache_aw_valid_o  (),
    .icache_aw_ready_i  (),
    .icache_ar_addr_o   (icache.ar_addr),
    .icache_ar_prot_o   (icache.ar_prot),
    .icache_ar_region_o (icache.ar_region),
    .icache_ar_len_o    (icache.ar_len),
    .icache_ar_size_o   (icache.ar_size),
    .icache_ar_burst_o  (icache.ar_burst),
    .icache_ar_lock_o   (icache.ar_lock),
    .icache_ar_cache_o  (icache.ar_cache),
    .icache_ar_qos_o    (icache.ar_qos),
    .icache_ar_id_o     (icache.ar_id),
    .icache_ar_user_o   (icache.ar_user),
    .icache_ar_valid_o  (),
    .icache_ar_ready_i  (),
    .icache_w_data_o    (icache.w_data),
    .icache_w_strb_o    (icache.w_strb),
    .icache_w_user_o    (icache.w_user),
    .icache_w_last_o    (icache.w_last),
    .icache_w_valid_o   (),
    .icache_w_ready_i   (),
    .icache_r_data_i    (icache.r_data),
    .icache_r_resp_i    (icache.r_resp),
    .icache_r_last_i    (icache.r_last),
    .icache_r_id_i      (icache.r_id),
    .icache_r_user_i    (icache.r_user),
    .icache_r_valid_i   (),
    .icache_r_ready_o   (),
    .icache_b_resp_i    (icache.b_resp),
    .icache_b_id_i      (icache.b_id),
    .icache_b_user_i    (icache.b_user),
    .icache_b_valid_i   (),
    .icache_b_ready_o   ()
  );
endmodule
